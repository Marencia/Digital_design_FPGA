library ieee;
use ieee.std_logic_1164.all;

entity contador_a is 
port ( clk, reset1: in std_logic;
			y: out std_logic_vector(3 downto 0)
		);
end contador_a;

architecture estructura of contador_a is
begin

process (clk)
	
	variable i: integer:=0;
	
begin

	if rising_edge(clk) then
		
		
		case i is
		
				when  0  =>	y<="0000";
				when  1  =>	y<="0001";
				when  2  =>	y<="0010";
				when  3  =>	y<="0011";
				when  4  =>	y<="0100";
				when  5  =>	y<="0101";
				when  6  =>	y<="0110";
				when  7  =>	y<="0111";
				when  8  =>	y<="1000";
				when  9  =>	y<="1001";
				when  10 =>	y<="1010";
				when  11 =>	y<="1011";
				when  12 =>	y<="1100";
				when  13 =>	y<="1101";
				when  14 =>	y<="1110";
				when  15 =>	y<="1111";
			
			when others =>	y<="ZZZZ";
					
		end case;
		i:=i+1;
		
	end if;
		
	if reset1 = '1' then
			i:=0;
	end if;
			
			
		
end process;
end estructura;