library ieee;
use ieee.std_logic_1164.all;

entity codificador_b is
port	(a: in std_logic_vector(7 downto 0);
		 y: out std_logic_vector (2 downto 0)
		 );
end codificador_b;

architecture estructura of  codificador_b is
begin

process (a)
begin

if a = "10000000" then 
	y<="111";
	
	elsif a = "01000000" then
		y<="110";
		
		elsif a = "00100000" then
			y<="101";
			
			elsif a = "00010000" then
				y<="100";
				
				elsif a = "00001000" then
					y<="011";
					
					elsif a = "00000100" then
						y<="010";
						
						elsif a = "00000010" then
							y<="001";
							
							elsif a = "00000001" then
								y<="000";
								
								else y<="ZZZ";
end if;		
end process;
end estructura;
